----------------------------------------------------------------------------------
-- Final Project
-- Processor
-- Baktash Ansari
-- Amir Reza Vishteh
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use std.textio.all;
use ieee.numeric_std.all;
use ieee.math_real.uniform;
use ieee.math_real.floor;


-- Explanation : The processor is a Black-Box component that generate random 16 bits virtual address 
-- from specific file.	

entity Processor is

port(
	

	index_file :  in integer;
	Output : out std_logic_vector(15 downto 0); -- virtual address
	read_bit : in std_logic
	
);

end Processor;

architecture Behavioral of Processor is



begin

--Generate random number from 0 to 199 . this number is the line number of file 
process is
	

	 variable rand_num : integer := 0;
    variable seed1 : positive;
    variable seed2 : positive;
    variable rand: real;   -- random real-number value in range 0 to 1.0  
    variable range_of_rand : real := 199.0;    -- the range of random values created will be 0 to +1000.
	 
	 
	 type addresses is array (0 to 199) of std_logic_vector(15 downto 0);
	 variable arry : addresses := (
		"1011001101010111",
		"1101110111010010",
		"1000000111001110",
		"0110111000000001",
		"1001001010100111",
		"1001011101000101",
		"0010100110100011",
		"1110010000111011",
		"0111011000000110",
		"0110110110110100",
		"1111011101011011",
		"0000110111011101",
		"0010110011110111",
		"0000100111101110",
		"0100111100110010",
		"1010011110010100",
		"1100111111010100",
		"1101010101100100",
		"1010001100100010",
		"1111100011000011",
		"1100011110100001",
		"0111101100101111",
		"1101111100011011",
		"1111111000011101",
		"1110111101011111",
		"1110100110111010",
		"0110010011001110",
		"0001000001010100",
		"1010111000100010",
		"1001110001001101",
		"1010100000101110",
		"0111100011010001",
		"1101001101010011",
		"1101111100100010",
		"0001110110110000",
		"0011001101111101",
		"1100001011110010",
		"1111001001000100",
		"0010010100100011",
		"1011000111001110",
		"0111011011011100",
		"0000001110101001",
		"0001011010110010",
		"0011011110110001",
		"1011100011011110",
		"0011111000010010",
		"1100101110011000",
		"0001010101010001",
		"1111100110010111",
		"0101001110110100",
		"0110100110001110",
		"0001111110001110",
		"0000111101110100",
		"1011111011001000",
		"1101011011100100",
		"1110001110110001",
		"0111101101110000",
		"1010010111100001",
		"0010110101110011",
		"0001101101000010",
		"1000101000100100",
		"0101101100010011",
		"1101111010000000",
		"0011110011110101",
		"1001111111101011",
		"1111010110111000",
		"1001101011011100",
		"1111111010100110",
		"1011000101010101",
		"1111010110011001",
		"0011101011011111",
		"1101010001110001",
		"1011001100100010",
		"1001000100100100",
		"1000111010110001",
		"1010110001000011",
		"0101010100101000",
		"0010101100110001",
		"0110101011010010",
		"0011000111010010",
		"1111100000100111",
		"0111010110101000",
		"1101101000111111",
		"0000010000000011",
		"0011111111100000",
		"1011011011101100",
		"1111011000110100",
		"0010011101100011",
		"0010011011011000",
		"1001000101111001",
		"0011010010001100",
		"0100011110110101",
		"0101100011010101",
		"1110110000001100",
		"0000100011111010",
		"1010101101111100",
		"1001010110000010",
		"1001010111100010",
		"0010011000010100",
		"1110111000011101",
		"0000110001010101",
		"0100100001001010",
		"1100111100101001",
		"1000011010111001",
		"1111101010101101",
		"1000000100000010",
		"1001100001000000",
		"1001001000110011",
		"0100100110111100",
		"0110000011110010",
		"1001101000000101",
		"1010101110010001",
		"0100110101001101",
		"0011000001000111",
		"1000010101101111",
		"0111101010111101",
		"1011011110001101",
		"0001011000010000",
		"0000010100001111",
		"1111000011011010",
		"1000010011110001",
		"1110001000000001",
		"1000000111000100",
		"0010101111000011",
		"0101111110001111",
		"1110101110111100",
		"1000101000010011",
		"1110000110010011",
		"0110111000001100",
		"0011110011001010",
		"1110011011010000",
		"0110101100010111",
		"1111110111001100",
		"1010111111001011",
		"1011111011111011",
		"1001010010001011",
		"0111111101111100",
		"1100011111101001",
		"1010010111100000",
		"0011101010000000",
		"1110011100000001",
		"1000001110000011",
		"0100000100000111",
		"0001100100111011",
		"1001111011101111",
		"0000100010100011",
		"1011010010001001",
		"0111111001111110",
		"0001111111011010",
		"0110001000101101",
		"1001011101110000",
		"1001101100110100",
		"1011000111001101",
		"0011011001101101",
		"0001011110111010",
		"0010101110011001",
		"1000111100000011",
		"0101100001010111",
		"1000100110101111",
		"0001101011000010",
		"1011011000101011",
		"0111001001001011",
		"1101110100101000",
		"0000001100011010",
		"1111110010110010",
		"1001111011001101",
		"1110100100001101",
		"1010010110011000",
		"1111001100101011",
		"1010001010101100",
		"1101100110011000",
		"1111001101110001",
		"0000000100010110",
		"1000010000001000",
		"1001011100011101",
		"0010110011110010",
		"1100111011001101",
		"1111000110001101",
		"0010010011111101",
		"1100001001110100",
		"1001011000100100",
		"1011110110101001",
		"1110110001101110",
		"1110010011100111",
		"0111100100111100",
		"1101100000100111",
		"0111000010110001",
		"0100000101100000",
		"0111100001110101",
		"0111010000011101",
		"1101100101011011",
		"0000011111110100",
		"0010111111000000",
		"0010011000111101",
		"0011000100111110",
		"1100110011001001",
		"1110000101110101",
		"0011010101001010",
		"1101110100001001",
		"0101100011000111"
);
  begin
    --uniform(seed1, seed2, rand);   -- generate random number
    --rand_num := integer(rand*range_of_rand);  -- rescale to 0..199, convert integer part 
    --wait for 10 ns;
	 if read_bit = '1' then
		Output <= arry(index_file);
	 end if;
	wait;
  end process;

end Behavioral;

